module example_combinational_1(input wire a, input wire b, output wire y,output wire x);
    assign y = a & b;
	 assign x = a ^ b;
endmodule




